output_buffer_inst : output_buffer PORT MAP (
		datain	 => datain_sig,
		oe	 => oe_sig,
		dataout	 => dataout_sig
	);
